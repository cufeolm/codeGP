`include "GUVM_test.sv"
`include"add_test.sv"
`include"bief_test.sv"
`include"child_test.sv"
`include"A_type_test.sv"
`include"subcc_test.sv"
`include"load_double_test.sv"
`include"arith_flag_test.sv"
`include"store_test.sv"
`include"mul_test.sv"
`include"arith_flag_amber_test.sv"


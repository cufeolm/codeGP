
// get_format switch case 
parameter REGOP_SWAP_MULT          = 3'b000;
parameter REGOP                    = 3'b001;
parameter TRANS_imm                = 3'b010;
parameter TRANS_reg                = 3'b011;
parameter MTRANS                   = 3'b100;
parameter BRANCH                   = 3'b101;
parameter CODTRANS                 = 3'b110;
parameter COREGOP_CORTRANS_SWI     = 3'b111;
function void verify_test(target_seq_item cmd_trans,GUVM_result_transaction res_trans);
	
endfunction
`include "riscy_pkg.sv"
`include "leon_seq_item.sv"
`include "GUVM_sequence.sv"
`include "child_sequence.sv"
`include "A_type_seq.sv"
`include"add_seq.sv"
`include"bief_seq.sv"
`include"subcc_seq.sv"
`include"load_double_seq.sv"
`include"arith_flag_seq.sv"
`include"store_seq.sv"
`include"mul_sequence.sv"


`include "leon_pkg.sv"
`include "GUVM_result_transaction.sv"
`include "GUVM_sequence_item.sv"
`include "target_sequence_item.sv"
`include "GUVM_sequence.sv"
`include "GUVM_driver.sv"
`include "GUVM_monitor.sv"
`include "GUVM_scoreboard.sv"
`include "GUVM_agent.sv"
`include "GUVM_env.sv"
`include "GUVM_test.sv"
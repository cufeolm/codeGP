`include "riscy_seq_item.sv"

// get_format switch case 
parameter U_type          = 7'b0110111;
parameter U_type1                    = 7'b0010111;
parameter J_type                = 7'b1101111;
parameter I_type                = 7'b1100111;
parameter I_type1                   = 7'b0000011;
parameter I_type_shift                   = 7'b0010011;
parameter I_type_fence                 = 7'b0001111;
parameter I_type_csr     = 7'b1110011;
parameter B_type                   = 7'b1100011;
parameter S_type                   = 7'b0100011;
parameter R_type                 = 7'b0110011;

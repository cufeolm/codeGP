`include "amber_seq_item.sv"
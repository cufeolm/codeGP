
// get_format switch case 
parameter CALL                            = 3'b00;
parameter SETHI_NOP_BRANCH                = 3'b01;
parameter Remaining_instructions          = 3'b10;
parameter Remaining_instructions1          = 3'b11;

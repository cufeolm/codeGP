// Da hayet7at feeh el interface elly hane5taro mn ay wa7ed mn rlfiles elly m3ana
`include "add.svh"
`include "test.svh"
`include "amber_pkg.sv"